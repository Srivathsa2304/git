module shrikanth;
  abcd 
  efgh
endmodule
