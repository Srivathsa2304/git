module shrikanth;
endmodule
